`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/04/2020 04:28:43 PM
// Design Name: 
// Module Name: Lab2A
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Lab2A(
    input [0:0] Read1,
    input [0:0] Read2,
    input [0:0] WriteReg,
    input [0:0] WriteData,
    input RegWrite,
    input clock,
    output [0:0] Data1,
    output [0:0] Data2
    );
endmodule
